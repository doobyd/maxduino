module maxduino
(
	input  wire		clk,
	input  wire		reset_n,
	input  wire		rxd,
	output wire		txd,
	output wire [21:0] gpio
);
	 
endmodule